VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
USEMINSPACING OBS OFF ;
CLEARANCEMEASURE EUCLIDEAN ;

UNITS
  DATABASE MICRONS 2000 ;
END UNITS

MANUFACTURINGGRID 0.0005 ;

PROPERTYDEFINITIONS
  LAYER LEF58_RIGHTWAYONGRIDONLY STRING ;
  LAYER LEF58_RECTONLY STRING ;
END PROPERTYDEFINITIONS

SITE coresite
    SIZE 0.045 BY 0.144 ;
    CLASS CORE ;
    SYMMETRY Y ;
END coresite
LAYER M0
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.024 ;
  OFFSET 0.0 ;
  WIDTH 0.014 ;
  MINWIDTH 0.014 ;
  AREA 0.000 ;
  SPACING 0.024 ENDOFLINE 0.024 WITHIN 0.001 ;
  SPACING 0.010 ;
  SPACINGTABLE  PARALLELRUNLENGTH
                0  
  WIDTH 0       0.010 ; 
  PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
  PROPERTY LEF58_RECTONLY " RECTONLY ; " ;
END M0
LAYER V0
  TYPE CUT ;
  WIDTH 0.012 ;
  SPACING 0.042 CENTERTOCENTER ;
END V0
LAYER M1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.030 ;
  OFFSET 0.0 ;
  WIDTH 0.015 ;
  MINWIDTH 0.015 ;
  AREA 0.000 ;
  SPACING 0.030 ENDOFLINE 0.030 WITHIN 0.001 ;
  SPACING 0.015 ;
  SPACINGTABLE  PARALLELRUNLENGTH
                0  
  WIDTH 0       0.015 ; 
  PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
  PROPERTY LEF58_RECTONLY " RECTONLY ; " ;
END M1
LAYER V1
  TYPE CUT ;
  WIDTH 0.014 ;
  SPACING 0.034 CENTERTOCENTER ;
END V1
LAYER M2
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.024 ;
  OFFSET 0.0 ;
  WIDTH 0.014 ;
  MINWIDTH 0.014 ;
  AREA 0.000 ;
  SPACING 0.024 ENDOFLINE 0.024 WITHIN 0.001 ;
  SPACING 0.010 ;
  SPACINGTABLE  PARALLELRUNLENGTH
                0  
  WIDTH 0       0.010 ; 
  PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
  PROPERTY LEF58_RECTONLY " RECTONLY ; " ;
END M2
LAYER V2
  TYPE CUT ;
  WIDTH 0.012 ;
  SPACING 0.034 CENTERTOCENTER ;
END V2
LAYER M3
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.024 ;
  OFFSET 0.0 ;
  WIDTH 0.014 ;
  MINWIDTH 0.014 ;
  AREA 0.000 ;
  SPACING 0.024 ENDOFLINE 0.024 WITHIN 0.001 ;
  SPACING 0.010 ;
  SPACINGTABLE  PARALLELRUNLENGTH
                0  
  WIDTH 0       0.010 ; 
  PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
  PROPERTY LEF58_RECTONLY " RECTONLY ; " ;
END M3
LAYER V3
  TYPE CUT ;
  WIDTH 0.012 ;
  SPACING 0.091 CENTERTOCENTER ;
END V3
LAYER M4
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.064 ;
  OFFSET 0.0 ;
  WIDTH 0.032 ;
  MINWIDTH 0.032 ;
  AREA 0.002 ;
  SPACING 0.064 ENDOFLINE 0.064 WITHIN 0.001 ;
  SPACING 0.032 ;
  SPACINGTABLE  PARALLELRUNLENGTH
                0  
  WIDTH 0       0.032 ; 
  PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
  PROPERTY LEF58_RECTONLY " RECTONLY ; " ;
END M4
LAYER V4
  TYPE CUT ;
  WIDTH 0.032 ;
  SPACING 0.091 CENTERTOCENTER ;
END V4
LAYER M5
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.064 ;
  OFFSET 0.0 ;
  WIDTH 0.032 ;
  MINWIDTH 0.032 ;
  AREA 0.002 ;
  SPACING 0.064 ENDOFLINE 0.064 WITHIN 0.001 ;
  SPACING 0.032 ;
  SPACINGTABLE  PARALLELRUNLENGTH
                0  
  WIDTH 0       0.032 ; 
  PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
  PROPERTY LEF58_RECTONLY " RECTONLY ; " ;
END M5
LAYER V5
  TYPE CUT ;
  WIDTH 0.032 ;
  SPACING 0.091 CENTERTOCENTER ;
END V5
LAYER M6
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.064 ;
  OFFSET 0.0 ;
  WIDTH 0.032 ;
  MINWIDTH 0.032 ;
  AREA 0.002 ;
  SPACING 0.064 ENDOFLINE 0.064 WITHIN 0.001 ;
  SPACING 0.032 ;
  SPACINGTABLE  PARALLELRUNLENGTH
                0  
  WIDTH 0       0.032 ; 
  PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
  PROPERTY LEF58_RECTONLY " RECTONLY ; " ;
END M6
LAYER V6
  TYPE CUT ;
  WIDTH 0.032 ;
  SPACING 0.091 CENTERTOCENTER ;
END V6
LAYER M7
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.064 ;
  OFFSET 0.0 ;
  WIDTH 0.032 ;
  MINWIDTH 0.032 ;
  AREA 0.002 ;
  SPACING 0.064 ENDOFLINE 0.064 WITHIN 0.001 ;
  SPACING 0.032 ;
  SPACINGTABLE  PARALLELRUNLENGTH
                0  
  WIDTH 0       0.032 ; 
  PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
  PROPERTY LEF58_RECTONLY " RECTONLY ; " ;
END M7
LAYER V7
  TYPE CUT ;
  WIDTH 0.032 ;
  SPACING 0.091 CENTERTOCENTER ;
END V7
LAYER M8
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.064 ;
  OFFSET 0.0 ;
  WIDTH 0.032 ;
  MINWIDTH 0.032 ;
  AREA 0.002 ;
  SPACING 0.064 ENDOFLINE 0.064 WITHIN 0.001 ;
  SPACING 0.032 ;
  SPACINGTABLE  PARALLELRUNLENGTH
                0  
  WIDTH 0       0.032 ; 
  PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
  PROPERTY LEF58_RECTONLY " RECTONLY ; " ;
END M8
LAYER V8
  TYPE CUT ;
  WIDTH 0.032 ;
  SPACING 0.091 CENTERTOCENTER ;
END V8
LAYER M9
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.064 ;
  OFFSET 0.0 ;
  WIDTH 0.032 ;
  MINWIDTH 0.032 ;
  AREA 0.002 ;
  SPACING 0.064 ENDOFLINE 0.064 WITHIN 0.001 ;
  SPACING 0.032 ;
  SPACINGTABLE  PARALLELRUNLENGTH
                0  
  WIDTH 0       0.032 ; 
  PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
  PROPERTY LEF58_RECTONLY " RECTONLY ; " ;
END M9
LAYER V9
  TYPE CUT ;
  WIDTH 0.032 ;
  SPACING 0.091 CENTERTOCENTER ;
END V9
LAYER M10
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.064 ;
  OFFSET 0.0 ;
  WIDTH 0.032 ;
  MINWIDTH 0.032 ;
  AREA 0.002 ;
  SPACING 0.064 ENDOFLINE 0.064 WITHIN 0.001 ;
  SPACING 0.032 ;
  SPACINGTABLE  PARALLELRUNLENGTH
                0  
  WIDTH 0       0.032 ; 
  PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
  PROPERTY LEF58_RECTONLY " RECTONLY ; " ;
END M10
LAYER V10
  TYPE CUT ;
  WIDTH 0.032 ;
  SPACING 0.091 CENTERTOCENTER ;
END V10
LAYER M11
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.064 ;
  OFFSET 0.0 ;
  WIDTH 0.032 ;
  MINWIDTH 0.032 ;
  AREA 0.002 ;
  SPACING 0.064 ENDOFLINE 0.064 WITHIN 0.001 ;
  SPACING 0.032 ;
  SPACINGTABLE  PARALLELRUNLENGTH
                0  
  WIDTH 0       0.032 ; 
  PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
  PROPERTY LEF58_RECTONLY " RECTONLY ; " ;
END M11
LAYER V11
  TYPE CUT ;
  WIDTH 0.032 ;
  SPACING 1.018 CENTERTOCENTER ;
END V11
LAYER M12
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.720 ;
  OFFSET 0.0 ;
  WIDTH 0.360 ;
  MINWIDTH 0.360 ;
  AREA 0.259 ;
  SPACING 0.720 ENDOFLINE 0.720 WITHIN 0.001 ;
  SPACING 0.360 ;
  SPACINGTABLE  PARALLELRUNLENGTH
                0  
  WIDTH 0       0.360 ; 
  PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
  PROPERTY LEF58_RECTONLY " RECTONLY ; " ;
END M12
LAYER V12
  TYPE CUT ;
  WIDTH 0.360 ;
  SPACING 1.018 CENTERTOCENTER ;
END V12
LAYER M13
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.720 ;
  OFFSET 0.0 ;
  WIDTH 0.360 ;
  MINWIDTH 0.360 ;
  AREA 0.259 ;
  SPACING 0.720 ENDOFLINE 0.720 WITHIN 0.001 ;
  SPACING 0.360 ;
  SPACINGTABLE  PARALLELRUNLENGTH
                0  
  WIDTH 0       0.360 ; 
  PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
  PROPERTY LEF58_RECTONLY " RECTONLY ; " ;
END M13
LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP
VIARULE V0_RULE GENERATE
  LAYER M0 ;
    ENCLOSURE 0.007 0.000 ;
  LAYER M1 ;
    ENCLOSURE 0.007 0.0004999999999999996 ;
  LAYER V0 ;
    RECT -0.007 -0.007 0.007 0.007 ;
    SPACING 0.042 BY 0.042 ;
END V0_RULE
VIARULE V1_RULE GENERATE
  LAYER M1 ;
    ENCLOSURE 0.007 0.0004999999999999996 ;
  LAYER M2 ;
    ENCLOSURE 0.007 0.000 ;
  LAYER V1 ;
    RECT -0.007 -0.007 0.007 0.007 ;
    SPACING 0.034 BY 0.034 ;
END V1_RULE
VIARULE V2_RULE GENERATE
  LAYER M2 ;
    ENCLOSURE 0.007 0.000 ;
  LAYER M3 ;
    ENCLOSURE 0.007 0.000 ;
  LAYER V2 ;
    RECT -0.007 -0.007 0.007 0.007 ;
    SPACING 0.034 BY 0.034 ;
END V2_RULE
VIARULE V3_RULE GENERATE
  LAYER M3 ;
    ENCLOSURE 0.007 0.000 ;
  LAYER M4 ;
    ENCLOSURE 0.007 0.009000000000000001 ;
  LAYER V3 ;
    RECT -0.007 -0.007 0.007 0.007 ;
    SPACING 0.091 BY 0.091 ;
END V3_RULE
VIARULE V4_RULE GENERATE
  LAYER M4 ;
    ENCLOSURE 0.007 0.000 ;
  LAYER M5 ;
    ENCLOSURE 0.007 0.000 ;
  LAYER V4 ;
    RECT -0.016 -0.016 0.016 0.016 ;
    SPACING 0.091 BY 0.091 ;
END V4_RULE
VIARULE V5_RULE GENERATE
  LAYER M5 ;
    ENCLOSURE 0.007 0.000 ;
  LAYER M6 ;
    ENCLOSURE 0.007 0.000 ;
  LAYER V5 ;
    RECT -0.016 -0.016 0.016 0.016 ;
    SPACING 0.091 BY 0.091 ;
END V5_RULE
VIARULE V6_RULE GENERATE
  LAYER M6 ;
    ENCLOSURE 0.007 0.000 ;
  LAYER M7 ;
    ENCLOSURE 0.007 0.000 ;
  LAYER V6 ;
    RECT -0.016 -0.016 0.016 0.016 ;
    SPACING 0.091 BY 0.091 ;
END V6_RULE
VIARULE V7_RULE GENERATE
  LAYER M7 ;
    ENCLOSURE 0.007 0.000 ;
  LAYER M8 ;
    ENCLOSURE 0.007 0.000 ;
  LAYER V7 ;
    RECT -0.016 -0.016 0.016 0.016 ;
    SPACING 0.091 BY 0.091 ;
END V7_RULE
VIARULE V8_RULE GENERATE
  LAYER M8 ;
    ENCLOSURE 0.007 0.000 ;
  LAYER M9 ;
    ENCLOSURE 0.007 0.000 ;
  LAYER V8 ;
    RECT -0.016 -0.016 0.016 0.016 ;
    SPACING 0.091 BY 0.091 ;
END V8_RULE
VIARULE V9_RULE GENERATE
  LAYER M9 ;
    ENCLOSURE 0.007 0.000 ;
  LAYER M10 ;
    ENCLOSURE 0.007 0.000 ;
  LAYER V9 ;
    RECT -0.016 -0.016 0.016 0.016 ;
    SPACING 0.091 BY 0.091 ;
END V9_RULE
VIARULE V10_RULE GENERATE
  LAYER M10 ;
    ENCLOSURE 0.007 0.000 ;
  LAYER M11 ;
    ENCLOSURE 0.007 0.000 ;
  LAYER V10 ;
    RECT -0.016 -0.016 0.016 0.016 ;
    SPACING 0.091 BY 0.091 ;
END V10_RULE
VIARULE V11_RULE GENERATE
  LAYER M11 ;
    ENCLOSURE 0.007 0.000 ;
  LAYER M12 ;
    ENCLOSURE 0.007 0.16399999999999998 ;
  LAYER V11 ;
    RECT -0.016 -0.016 0.016 0.016 ;
    SPACING 1.018 BY 1.018 ;
END V11_RULE
VIARULE V12_RULE GENERATE
  LAYER M12 ;
    ENCLOSURE 0.007 0.000 ;
  LAYER M13 ;
    ENCLOSURE 0.007 0.000 ;
  LAYER V12 ;
    RECT -0.180 -0.180 0.180 0.180 ;
    SPACING 1.018 BY 1.018 ;
END V12_RULE
VIA V0_HV DEFAULT
  LAYER M0 ;
  RECT -0.014 -0.007 0.014 0.007 ;
  LAYER V0 ;
  RECT -0.007 -0.007 0.007 0.007 ;
  LAYER M1 ;
  RECT -0.007 -0.014 0.007 0.014 ;
END V0_HV
VIA V1_VH DEFAULT
  LAYER M1 ;
  RECT -0.007 -0.014 0.007 0.014 ;
  LAYER V1 ;
  RECT -0.007 -0.007 0.007 0.007 ;
  LAYER M2 ;
  RECT -0.014 -0.007 0.014 0.007 ;
END V1_VH
VIA V2_HV DEFAULT
  LAYER M2 ;
  RECT -0.014 -0.007 0.014 0.007 ;
  LAYER V2 ;
  RECT -0.007 -0.007 0.007 0.007 ;
  LAYER M3 ;
  RECT -0.007 -0.014 0.007 0.014 ;
END V2_HV
VIA V3_VH DEFAULT
  LAYER M3 ;
  RECT -0.007 -0.014 0.007 0.014 ;
  LAYER V3 ;
  RECT -0.007 -0.007 0.007 0.007 ;
  LAYER M4 ;
  RECT -0.014 -0.016 0.014 0.016 ;
END V3_VH
VIA V4_HV DEFAULT
  LAYER M4 ;
  RECT -0.023 -0.016 0.023 0.016 ;
  LAYER V4 ;
  RECT -0.016 -0.016 0.016 0.016 ;
  LAYER M5 ;
  RECT -0.016 -0.023 0.016 0.023 ;
END V4_HV
VIA V5_VH DEFAULT
  LAYER M5 ;
  RECT -0.016 -0.023 0.016 0.023 ;
  LAYER V5 ;
  RECT -0.016 -0.016 0.016 0.016 ;
  LAYER M6 ;
  RECT -0.023 -0.016 0.023 0.016 ;
END V5_VH
VIA V6_HV DEFAULT
  LAYER M6 ;
  RECT -0.023 -0.016 0.023 0.016 ;
  LAYER V6 ;
  RECT -0.016 -0.016 0.016 0.016 ;
  LAYER M7 ;
  RECT -0.016 -0.023 0.016 0.023 ;
END V6_HV
VIA V7_VH DEFAULT
  LAYER M7 ;
  RECT -0.016 -0.023 0.016 0.023 ;
  LAYER V7 ;
  RECT -0.016 -0.016 0.016 0.016 ;
  LAYER M8 ;
  RECT -0.023 -0.016 0.023 0.016 ;
END V7_VH
VIA V8_HV DEFAULT
  LAYER M8 ;
  RECT -0.023 -0.016 0.023 0.016 ;
  LAYER V8 ;
  RECT -0.016 -0.016 0.016 0.016 ;
  LAYER M9 ;
  RECT -0.016 -0.023 0.016 0.023 ;
END V8_HV
VIA V9_VH DEFAULT
  LAYER M9 ;
  RECT -0.016 -0.023 0.016 0.023 ;
  LAYER V9 ;
  RECT -0.016 -0.016 0.016 0.016 ;
  LAYER M10 ;
  RECT -0.023 -0.016 0.023 0.016 ;
END V9_VH
VIA V10_HV DEFAULT
  LAYER M10 ;
  RECT -0.023 -0.016 0.023 0.016 ;
  LAYER V10 ;
  RECT -0.016 -0.016 0.016 0.016 ;
  LAYER M11 ;
  RECT -0.016 -0.023 0.016 0.023 ;
END V10_HV
VIA V11_VH DEFAULT
  LAYER M11 ;
  RECT -0.016 -0.023 0.016 0.023 ;
  LAYER V11 ;
  RECT -0.016 -0.016 0.016 0.016 ;
  LAYER M12 ;
  RECT -0.023 -0.180 0.023 0.180 ;
END V11_VH
VIA V12_HV DEFAULT
  LAYER M12 ;
  RECT -0.187 -0.180 0.187 0.180 ;
  LAYER V12 ;
  RECT -0.180 -0.180 0.180 0.180 ;
  LAYER M13 ;
  RECT -0.180 -0.187 0.180 0.187 ;
END V12_HV
END LIBRARY
